`timescale 1ns / 1ps

// Encodes parallel HDMI commands for output
//
// The commands are presented over an AXI4-Stream slave interface. The input
// should likely have a FIFO to buffer commands, as this module will
// unconditionally request one command every cycle. The output should also be
// connected directly to the output pads, as this module takes care of
// generating the differential signals.
//
// Ports:
// * clk_px: Pixel clock. Should be 25.175MHz.
// * clk_5px: Clock that runs at 5x the pixel clock rate. It must be in phase
//   with `clk_px`. So for example, it could be generated by the same MMCM as
//   `clk_px`.
// * resetn_async: Active-low asynchronous reset. This can be tied to the
//   `locked` output of the clock generator.
// * commands: Interface on which HDMI commands are consumed. The LSB is the
//   first bit to be serialized. Bits [9:0] are the command for channel 0,
//   [19:10] for channel 1, and [29:20] for channel 2.
// * hdmi_pulse: Channel C for the HDMI output
// * hdmi_data: Serialized data for each channel. Bit 0 is for channel 0, bit 1
//   for channel 1, and bit 2 for channel 2.
module top(
    input clk_px,
    input clk_5px,
    input resetn_async,

    input [31:0] commands_tdata,
    input commands_tvalid,
    output commands_tready,

    output hdmi_pulse_p,
    output hdmi_pulse_n,
    output [2:0] hdmi_data_p,
    output [2:0] hdmi_data_n
);

// HDMI command corresponding to no active video and no synchronization signal
localparam HDMI_CMD_NOOP = 10'b1101010100;

// The input reset signal is asynchronous. However, the serializer requires that
// the reset be synchronous, and it's just good practice to have it. So,
// synchronize.
wire resetn;
wire reset;
reset_controller #(
    .NUM_STAGES(2)
) reset_controller (
    .clk(clk_px),
    .resetn_async(resetn_async),
    .resetn(resetn),
    .reset(reset)
);

// We consume one command every cycle, so we're always ready
assign commands_tready = 1'b1;

// If we're in reset, disable the output pulses and send noops. Otherwise, send
// the pulses and the input data. If the input data is not valid, just send
// noops. Put them in registers so we don't have a combinatorial path leading up
// to the serializers.
reg [9:0] hdmi_pulse;
reg [29:0] hdmi_data;
always @(posedge clk_px) begin
    if (resetn == 1'b0) begin
        hdmi_pulse <= 10'b0000000000;
        hdmi_data <= {3{HDMI_CMD_NOOP}};
    end else begin
        hdmi_pulse <= 10'b1111100000;
        if (commands_tvalid == 1'b1) begin
            hdmi_data <= commands_tdata[29:0];
        end else begin
            hdmi_data <= {3{HDMI_CMD_NOOP}};
        end
    end
end

// Serialize the clock pulse...
serializer pulse_ser(
    .clk_px(clk_px),
    .clk_5px(clk_5px),
    .reset(reset),
    .cmd(hdmi_pulse),
    .cmd_p(hdmi_pulse_p),
    .cmd_n(hdmi_pulse_n)
);
// ... as well as each of the channels
generate
for (genvar i = 0; i < 3; i = i + 1) begin
    serializer data_ser(
        .clk_px(clk_px),
        .clk_5px(clk_5px),
        .reset(reset),
        .cmd(hdmi_data[10*i+9:10*i]),
        .cmd_p(hdmi_data_p[i]),
        .cmd_n(hdmi_data_n[i])
    );
end
endgenerate

endmodule
