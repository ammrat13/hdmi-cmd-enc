`timescale 1ns / 1ps

// Serializer for a single TMDS channel
//
// We receive 10 bits of data in parallel for each channel. The job of this
// module is to serially put those bits on the output pin. To do this, it uses
// the OSERDES2 modules built in to each output buffer. It runs them in DDR
// mode, which means this module only needs a clock at 5x the pixel clock
// instead of 10x.
//
// Additionally, this module converts the logic signal inside the FPGA to a
// differential signal for output. The output ports with the serialized command
// should therefore be connected directly to the pads.
//
// See: UG471
//
// Ports:
// * clk_px: Pixel clock. Should be 25.175MHz.
// * clk_5px: Clock that runs at 5x the pixel clock rate. It must be in phase
//   with `clk_px`. So for example, it could be generated by the same MMCM as
//   `clk_px`.
// * reset: Synchronous active-high reset
// * cmd: The command to serialize. The LSB is the first bit serialized.
// * cmd_p: The serialized command's positive end of the differential pair
// * cmd_n: The serialized command's negative end of the differential pair
module serializer(
    input clk_px,
    input clk_5px,
    input reset,

    input [9:0] cmd,
    output cmd_p,
    output cmd_n
);

// This wire holds the output of the serializer while it's still a logic-level
// and not yet differential
wire cmd_s;

// Convert the logic-level serialized output to a differential signal
//
// See: UG471 Pg. 45
// See: https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/OBUFDS
OBUFDS #(
   .IOSTANDARD("TMDS_33"),
   .SLEW("SLOW")
) obuf (
   .O(cmd_p),
   .OB(cmd_n),
   .I(cmd_s)
);

// Setup the OSERDES2 modules for 10-bit serialization. We need two modules -
// one in master mode and one in slave mode. We don't use the tristate output
// functionality, so we tie the clock enable for it low and set the relevant
// parameters to silence warnings.
//
// See: UG471 Pg. 161
wire shift1;
wire shift2;
OSERDESE2 #(
   .DATA_RATE_OQ("DDR"),
   .DATA_WIDTH(10),
   .DATA_RATE_TQ("SDR"),
   .TRISTATE_WIDTH(1),
   .SERDES_MODE("MASTER")
) ser_master (
   .RST(reset),
   .CLK(clk_5px),
   .CLKDIV(clk_px),
   .OCE(1'b1),
   .TCE(1'b0),
   .D1(cmd[0]),
   .D2(cmd[1]),
   .D3(cmd[2]),
   .D4(cmd[3]),
   .D5(cmd[4]),
   .D6(cmd[5]),
   .D7(cmd[6]),
   .D8(cmd[7]),
   .OQ(cmd_s),
   .SHIFTIN1(shift1),
   .SHIFTIN2(shift2)
);
OSERDESE2 #(
   .DATA_RATE_OQ("DDR"),
   .DATA_WIDTH(10),
   .DATA_RATE_TQ("SDR"),
   .TRISTATE_WIDTH(1),
   .SERDES_MODE("SLAVE")
) ser_slave (
   .RST(reset),
   .CLK(clk_5px),
   .CLKDIV(clk_px),
   .OCE(1'b1),
   .TCE(1'b0),
   .D1(1'b0),
   .D2(1'b0),
   .D3(cmd[8]),
   .D4(cmd[9]),
   .D5(1'b0),
   .D6(1'b0),
   .D7(1'b0),
   .D8(1'b0),
   .SHIFTOUT1(shift1),
   .SHIFTOUT2(shift2)
);

endmodule
